------------------------------------------------------------------------------
----                                                                      ----
----  Dual Port RAM that maps to a Xilinx BRAM                            ----
----                                                                      ----
----  http://www.opencores.org/                                           ----
----                                                                      ----
----  Description:                                                        ----
----  This is a program+data memory for the ZPU. It maps to a Xilinx BRAM ----
----                                                                      ----
----  To Do:                                                              ----
----  -                                                                   ----
----                                                                      ----
----  Author:                                                             ----
----    - �yvind Harboe, oyvind.harboe zylin.com                          ----
----    - Salvador E. Tropea, salvador inti.gob.ar                        ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Copyright (c) 2008 �yvind Harboe <oyvind.harboe zylin.com>           ----
---- Copyright (c) 2008 Salvador E. Tropea <salvador inti.gob.ar>         ----
---- Copyright (c) 2008 Instituto Nacional de Tecnolog�a Industrial       ----
----                                                                      ----
---- Distributed under the BSD license                                    ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Design unit:      DualPortRAM(Xilinx) (Entity and architecture)      ----
---- File name:        rom.in.vhdl (template used)                        ----
---- Note:             None                                               ----
---- Limitations:      None known                                         ----
---- Errors:           None known                                         ----
---- Library:          work                                               ----
---- Dependencies:     IEEE.std_logic_1164                                ----
----                   IEEE.numeric_std                                   ----
---- Target FPGA:      Spartan 3 (XC3S1500-4-FG456)                       ----
---- Language:         VHDL                                               ----
---- Wishbone:         No                                                 ----
---- Synthesis tools:  Xilinx Release 9.2.03i - xst J.39                  ----
---- Simulation tools: GHDL [Sokcho edition] (0.2x)                       ----
---- Text editor:      SETEdit 0.5.x                                      ----
----                                                                      ----
------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DualPortRAM is
   generic(
      WORD_SIZE    : integer:=32;  -- Word Size 16/32
      BYTE_BITS    : integer:=2;   -- Bits used to address bytes
      BRAM_W       : integer:=15); -- Address Width
   port(
      clk_i     : in  std_logic;
      -- Port A
      a_we_i    : in  std_logic;
      a_addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      a_write_i : in  unsigned(WORD_SIZE-1 downto 0);
      a_read_o  : out unsigned(WORD_SIZE-1 downto 0);
      -- Port B
      b_we_i    : in  std_logic;
      b_addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      b_write_i : in  unsigned(WORD_SIZE-1 downto 0);
      b_read_o  : out unsigned(WORD_SIZE-1 downto 0));
end entity DualPortRAM;

architecture Xilinx of DualPortRAM is
   type ram_type is array(natural range 0 to ((2**BRAM_W)/4)-1) of unsigned(WORD_SIZE-1 downto 0);

   shared variable ram : ram_type:=
(
0 => x"0b0b0b0b",
1 => x"82700b0b",
2 => x"80d3e40c",
3 => x"3a0b0b80",
4 => x"cbba0400",
5 => x"00000000",
6 => x"00000000",
7 => x"00000000",
8 => x"0b0b0b89",
9 => x"90040000",
10 => x"00000000",
11 => x"00000000",
12 => x"00000000",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c4040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"020d0406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04000000",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80d3",
162 => x"80738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88aa0400",
166 => x"00000000",
167 => x"00000000",
168 => x"0b0b0b88",
169 => x"f8040000",
170 => x"00000000",
171 => x"00000000",
172 => x"00000000",
173 => x"00000000",
174 => x"00000000",
175 => x"00000000",
176 => x"0b0b0b88",
177 => x"e0040000",
178 => x"00000000",
179 => x"00000000",
180 => x"00000000",
181 => x"00000000",
182 => x"00000000",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07515151",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075151",
199 => x"51040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80d3e00c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"020d0400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"83863f80",
257 => x"cacd3f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51047381",
267 => x"ff067383",
268 => x"06098105",
269 => x"83051010",
270 => x"102b0772",
271 => x"fc060c51",
272 => x"51043c04",
273 => x"72728072",
274 => x"8106ff05",
275 => x"09720605",
276 => x"71105272",
277 => x"0a100a53",
278 => x"72ed3851",
279 => x"51535104",
280 => x"b008b408",
281 => x"b8087575",
282 => x"8ecf2d50",
283 => x"50b00856",
284 => x"b80cb40c",
285 => x"b00c5104",
286 => x"b008b408",
287 => x"b8087575",
288 => x"8d9d2d50",
289 => x"50b00856",
290 => x"b80cb40c",
291 => x"b00c5104",
292 => x"b008b408",
293 => x"b80880cc",
294 => x"852db80c",
295 => x"b40cb00c",
296 => x"04fe3d0d",
297 => x"0b0b80e3",
298 => x"cc085384",
299 => x"13087088",
300 => x"2a708106",
301 => x"51525270",
302 => x"802ef038",
303 => x"7181ff06",
304 => x"b00c843d",
305 => x"0d04ff3d",
306 => x"0d0b0b80",
307 => x"e3cc0852",
308 => x"71087088",
309 => x"2a813270",
310 => x"81065151",
311 => x"5170f138",
312 => x"73720c83",
313 => x"3d0d0480",
314 => x"d3e00880",
315 => x"2ea43880",
316 => x"d3e40882",
317 => x"2ebd3883",
318 => x"80800b0b",
319 => x"0b80e3cc",
320 => x"0c82a080",
321 => x"0b80e3d0",
322 => x"0c829080",
323 => x"0b80e3d4",
324 => x"0c04f880",
325 => x"8080a40b",
326 => x"0b0b80e3",
327 => x"cc0cf880",
328 => x"8082800b",
329 => x"80e3d00c",
330 => x"f8808084",
331 => x"800b80e3",
332 => x"d40c0480",
333 => x"c0a8808c",
334 => x"0b0b0b80",
335 => x"e3cc0c80",
336 => x"c0a88094",
337 => x"0b80e3d0",
338 => x"0c80d390",
339 => x"0b80e3d4",
340 => x"0c04ff3d",
341 => x"0d80e3d8",
342 => x"335170a7",
343 => x"3880d3ec",
344 => x"08700852",
345 => x"5270802e",
346 => x"94388412",
347 => x"80d3ec0c",
348 => x"702d80d3",
349 => x"ec087008",
350 => x"525270ee",
351 => x"38810b80",
352 => x"e3d83483",
353 => x"3d0d0404",
354 => x"803d0d0b",
355 => x"0b80e3c8",
356 => x"08802e8e",
357 => x"380b0b0b",
358 => x"0b800b80",
359 => x"2e098106",
360 => x"8538823d",
361 => x"0d040b0b",
362 => x"80e3c851",
363 => x"0b0b0bf4",
364 => x"cf3f823d",
365 => x"0d0404fd",
366 => x"3d0d8170",
367 => x"54547280",
368 => x"c0a88084",
369 => x"0c80c0a8",
370 => x"80840870",
371 => x"822a8106",
372 => x"70307072",
373 => x"07700970",
374 => x"9f2c7906",
375 => x"781081fe",
376 => x"06595951",
377 => x"51535152",
378 => x"72833881",
379 => x"5373cf38",
380 => x"853d0d04",
381 => x"ff3d0d80",
382 => x"c0a88084",
383 => x"5282d480",
384 => x"80720c80",
385 => x"c0a88088",
386 => x"51f883ff",
387 => x"ff710c85",
388 => x"a8808072",
389 => x"0cff710c",
390 => x"833d0d04",
391 => x"fc3d0d80",
392 => x"d3945186",
393 => x"da3f80d3",
394 => x"a05186d3",
395 => x"3f80d3b0",
396 => x"5186cc3f",
397 => x"81705555",
398 => x"7380c0a8",
399 => x"80840c80",
400 => x"c0a88084",
401 => x"0870822a",
402 => x"81067030",
403 => x"70720770",
404 => x"09709f2c",
405 => x"7a067910",
406 => x"81fe065a",
407 => x"5a515154",
408 => x"51537383",
409 => x"38815474",
410 => x"cf3882d4",
411 => x"80800b80",
412 => x"c0a88084",
413 => x"0cf883ff",
414 => x"ff0b80c0",
415 => x"a880880c",
416 => x"85a88080",
417 => x"0b80c0a8",
418 => x"80840cff",
419 => x"0b80c0a8",
420 => x"80880c80",
421 => x"d3c05185",
422 => x"e63f83fd",
423 => x"3fbc0802",
424 => x"bc0cf93d",
425 => x"0d800bbc",
426 => x"08fc050c",
427 => x"bc088805",
428 => x"088025ab",
429 => x"38bc0888",
430 => x"050830bc",
431 => x"0888050c",
432 => x"800bbc08",
433 => x"f4050cbc",
434 => x"08fc0508",
435 => x"8838810b",
436 => x"bc08f405",
437 => x"0cbc08f4",
438 => x"0508bc08",
439 => x"fc050cbc",
440 => x"088c0508",
441 => x"8025ab38",
442 => x"bc088c05",
443 => x"0830bc08",
444 => x"8c050c80",
445 => x"0bbc08f0",
446 => x"050cbc08",
447 => x"fc050888",
448 => x"38810bbc",
449 => x"08f0050c",
450 => x"bc08f005",
451 => x"08bc08fc",
452 => x"050c8053",
453 => x"bc088c05",
454 => x"0852bc08",
455 => x"88050851",
456 => x"81a73fb0",
457 => x"0870bc08",
458 => x"f8050c54",
459 => x"bc08fc05",
460 => x"08802e8c",
461 => x"38bc08f8",
462 => x"050830bc",
463 => x"08f8050c",
464 => x"bc08f805",
465 => x"0870b00c",
466 => x"54893d0d",
467 => x"bc0c04bc",
468 => x"0802bc0c",
469 => x"fb3d0d80",
470 => x"0bbc08fc",
471 => x"050cbc08",
472 => x"88050880",
473 => x"259338bc",
474 => x"08880508",
475 => x"30bc0888",
476 => x"050c810b",
477 => x"bc08fc05",
478 => x"0cbc088c",
479 => x"05088025",
480 => x"8c38bc08",
481 => x"8c050830",
482 => x"bc088c05",
483 => x"0c8153bc",
484 => x"088c0508",
485 => x"52bc0888",
486 => x"050851ad",
487 => x"3fb00870",
488 => x"bc08f805",
489 => x"0c54bc08",
490 => x"fc050880",
491 => x"2e8c38bc",
492 => x"08f80508",
493 => x"30bc08f8",
494 => x"050cbc08",
495 => x"f8050870",
496 => x"b00c5487",
497 => x"3d0dbc0c",
498 => x"04bc0802",
499 => x"bc0cfd3d",
500 => x"0d810bbc",
501 => x"08fc050c",
502 => x"800bbc08",
503 => x"f8050cbc",
504 => x"088c0508",
505 => x"bc088805",
506 => x"0827ac38",
507 => x"bc08fc05",
508 => x"08802ea3",
509 => x"38800bbc",
510 => x"088c0508",
511 => x"249938bc",
512 => x"088c0508",
513 => x"10bc088c",
514 => x"050cbc08",
515 => x"fc050810",
516 => x"bc08fc05",
517 => x"0cc939bc",
518 => x"08fc0508",
519 => x"802e80c9",
520 => x"38bc088c",
521 => x"0508bc08",
522 => x"88050826",
523 => x"a138bc08",
524 => x"880508bc",
525 => x"088c0508",
526 => x"31bc0888",
527 => x"050cbc08",
528 => x"f80508bc",
529 => x"08fc0508",
530 => x"07bc08f8",
531 => x"050cbc08",
532 => x"fc050881",
533 => x"2abc08fc",
534 => x"050cbc08",
535 => x"8c050881",
536 => x"2abc088c",
537 => x"050cffaf",
538 => x"39bc0890",
539 => x"0508802e",
540 => x"8f38bc08",
541 => x"88050870",
542 => x"bc08f405",
543 => x"0c518d39",
544 => x"bc08f805",
545 => x"0870bc08",
546 => x"f4050c51",
547 => x"bc08f405",
548 => x"08b00c85",
549 => x"3d0dbc0c",
550 => x"04803d0d",
551 => x"865184e7",
552 => x"3f8151ba",
553 => x"dd3ffc3d",
554 => x"0d767079",
555 => x"7b555555",
556 => x"558f7227",
557 => x"8c387275",
558 => x"07830651",
559 => x"70802ea7",
560 => x"38ff1252",
561 => x"71ff2e98",
562 => x"38727081",
563 => x"05543374",
564 => x"70810556",
565 => x"34ff1252",
566 => x"71ff2e09",
567 => x"8106ea38",
568 => x"74b00c86",
569 => x"3d0d0474",
570 => x"51727084",
571 => x"05540871",
572 => x"70840553",
573 => x"0c727084",
574 => x"05540871",
575 => x"70840553",
576 => x"0c727084",
577 => x"05540871",
578 => x"70840553",
579 => x"0c727084",
580 => x"05540871",
581 => x"70840553",
582 => x"0cf01252",
583 => x"718f26c9",
584 => x"38837227",
585 => x"95387270",
586 => x"84055408",
587 => x"71708405",
588 => x"530cfc12",
589 => x"52718326",
590 => x"ed387054",
591 => x"ff8339f7",
592 => x"3d0d7c70",
593 => x"525384bd",
594 => x"3f7254b0",
595 => x"085580d3",
596 => x"cc568157",
597 => x"b0088105",
598 => x"5a8b3de4",
599 => x"11595382",
600 => x"59f41352",
601 => x"7b881108",
602 => x"525384f8",
603 => x"3fb00830",
604 => x"70b00807",
605 => x"9f2c8a07",
606 => x"b00c538b",
607 => x"3d0d04ff",
608 => x"3d0d7352",
609 => x"80d3f008",
610 => x"51ffb43f",
611 => x"833d0d04",
612 => x"fd3d0d75",
613 => x"5384d813",
614 => x"08802e8a",
615 => x"38805372",
616 => x"b00c853d",
617 => x"0d048180",
618 => x"5272518a",
619 => x"9d3fb008",
620 => x"84d8140c",
621 => x"ff53b008",
622 => x"802ee438",
623 => x"b008549f",
624 => x"53807470",
625 => x"8405560c",
626 => x"ff135380",
627 => x"7324ce38",
628 => x"80747084",
629 => x"05560cff",
630 => x"13537280",
631 => x"25e338ff",
632 => x"bc39fd3d",
633 => x"0d757755",
634 => x"539f7427",
635 => x"8d389673",
636 => x"0cff5271",
637 => x"b00c853d",
638 => x"0d0484d8",
639 => x"13085271",
640 => x"802e9338",
641 => x"73101012",
642 => x"70087972",
643 => x"0c515271",
644 => x"b00c853d",
645 => x"0d047251",
646 => x"fef63fff",
647 => x"52b008d3",
648 => x"3884d813",
649 => x"08741010",
650 => x"1170087a",
651 => x"720c5151",
652 => x"52dd39f9",
653 => x"3d0d797b",
654 => x"5856769f",
655 => x"2680e838",
656 => x"84d81608",
657 => x"5473802e",
658 => x"aa387610",
659 => x"10147008",
660 => x"55557380",
661 => x"2eba3880",
662 => x"5873812e",
663 => x"8f3873ff",
664 => x"2ea33880",
665 => x"750c7651",
666 => x"732d8058",
667 => x"77b00c89",
668 => x"3d0d0475",
669 => x"51fe993f",
670 => x"ff58b008",
671 => x"ef3884d8",
672 => x"160854c6",
673 => x"3996760c",
674 => x"810bb00c",
675 => x"893d0d04",
676 => x"755181ed",
677 => x"3f7653b0",
678 => x"08527551",
679 => x"81ad3fb0",
680 => x"08b00c89",
681 => x"3d0d0496",
682 => x"760cff0b",
683 => x"b00c893d",
684 => x"0d04fc3d",
685 => x"0d767856",
686 => x"53ff5474",
687 => x"9f26b138",
688 => x"84d81308",
689 => x"5271802e",
690 => x"ae387410",
691 => x"10127008",
692 => x"53538154",
693 => x"71802e98",
694 => x"38825471",
695 => x"ff2e9138",
696 => x"83547181",
697 => x"2e8a3880",
698 => x"730c7451",
699 => x"712d8054",
700 => x"73b00c86",
701 => x"3d0d0472",
702 => x"51fd953f",
703 => x"b008f138",
704 => x"84d81308",
705 => x"52c439ff",
706 => x"3d0d7352",
707 => x"80d3f008",
708 => x"51fea03f",
709 => x"833d0d04",
710 => x"fe3d0d75",
711 => x"53745280",
712 => x"d3f00851",
713 => x"fdbc3f84",
714 => x"3d0d0480",
715 => x"3d0d80d3",
716 => x"f00851fc",
717 => x"db3f823d",
718 => x"0d04ff3d",
719 => x"0d735280",
720 => x"d3f00851",
721 => x"feec3f83",
722 => x"3d0d04fc",
723 => x"3d0d800b",
724 => x"80e3e40c",
725 => x"78527751",
726 => x"b49a3fb0",
727 => x"0854b008",
728 => x"ff2e8838",
729 => x"73b00c86",
730 => x"3d0d0480",
731 => x"e3e40855",
732 => x"74802ef0",
733 => x"38767571",
734 => x"0c5373b0",
735 => x"0c863d0d",
736 => x"04b3ec3f",
737 => x"04fd3d0d",
738 => x"75707183",
739 => x"06535552",
740 => x"70b83871",
741 => x"70087009",
742 => x"f7fbfdff",
743 => x"120670f8",
744 => x"84828180",
745 => x"06515152",
746 => x"53709d38",
747 => x"84137008",
748 => x"7009f7fb",
749 => x"fdff1206",
750 => x"70f88482",
751 => x"81800651",
752 => x"51525370",
753 => x"802ee538",
754 => x"72527133",
755 => x"5170802e",
756 => x"8a388112",
757 => x"70335252",
758 => x"70f83871",
759 => x"7431b00c",
760 => x"853d0d04",
761 => x"f23d0d60",
762 => x"62881108",
763 => x"7057575f",
764 => x"5a74802e",
765 => x"818f388c",
766 => x"1a227083",
767 => x"2a813270",
768 => x"81065155",
769 => x"58738638",
770 => x"901a0891",
771 => x"3879519c",
772 => x"cc3fff54",
773 => x"b00880ed",
774 => x"388c1a22",
775 => x"587d0857",
776 => x"807883ff",
777 => x"ff067081",
778 => x"2a708106",
779 => x"51565755",
780 => x"73752e80",
781 => x"d7387490",
782 => x"38760884",
783 => x"18088819",
784 => x"59565974",
785 => x"802ef238",
786 => x"74548880",
787 => x"75278438",
788 => x"88805473",
789 => x"5378529c",
790 => x"1a0851a4",
791 => x"1a085473",
792 => x"2d800bb0",
793 => x"082582e6",
794 => x"38b00819",
795 => x"75b00831",
796 => x"7f880508",
797 => x"b0083170",
798 => x"6188050c",
799 => x"56565973",
800 => x"ffb43880",
801 => x"5473b00c",
802 => x"903d0d04",
803 => x"75813270",
804 => x"81067641",
805 => x"51547380",
806 => x"2e81c138",
807 => x"74903876",
808 => x"08841808",
809 => x"88195956",
810 => x"5974802e",
811 => x"f238881a",
812 => x"087883ff",
813 => x"ff067089",
814 => x"2a708106",
815 => x"51565956",
816 => x"73802e82",
817 => x"fa387575",
818 => x"278d3877",
819 => x"872a7081",
820 => x"06515473",
821 => x"82b53874",
822 => x"76278338",
823 => x"74567553",
824 => x"78527908",
825 => x"5190f83f",
826 => x"881a0876",
827 => x"31881b0c",
828 => x"7908167a",
829 => x"0c745675",
830 => x"19757731",
831 => x"7f880508",
832 => x"78317061",
833 => x"88050c56",
834 => x"56597380",
835 => x"2efef438",
836 => x"8c1a2258",
837 => x"ff863977",
838 => x"78547953",
839 => x"7b525690",
840 => x"be3f881a",
841 => x"08783188",
842 => x"1b0c7908",
843 => x"187a0c7c",
844 => x"76315d7c",
845 => x"8e387951",
846 => x"9c863fb0",
847 => x"08818f38",
848 => x"b0085f75",
849 => x"19757731",
850 => x"7f880508",
851 => x"78317061",
852 => x"88050c56",
853 => x"56597380",
854 => x"2efea838",
855 => x"74818338",
856 => x"76088418",
857 => x"08881959",
858 => x"56597480",
859 => x"2ef23874",
860 => x"538a5278",
861 => x"518ec93f",
862 => x"b0087931",
863 => x"81055db0",
864 => x"08843881",
865 => x"155d815f",
866 => x"7c58747d",
867 => x"27833874",
868 => x"58941a08",
869 => x"881b0811",
870 => x"575c807a",
871 => x"085c5490",
872 => x"1a087b27",
873 => x"83388154",
874 => x"75782584",
875 => x"3873ba38",
876 => x"7b7824fe",
877 => x"e2387b53",
878 => x"78529c1a",
879 => x"0851a41a",
880 => x"0854732d",
881 => x"b00856b0",
882 => x"088024fe",
883 => x"e2388c1a",
884 => x"2280c007",
885 => x"54738c1b",
886 => x"23ff5473",
887 => x"b00c903d",
888 => x"0d047eff",
889 => x"a338ff87",
890 => x"39755378",
891 => x"527a518e",
892 => x"ee3f7908",
893 => x"167a0c79",
894 => x"519ac53f",
895 => x"b008cf38",
896 => x"7c76315d",
897 => x"7cfebc38",
898 => x"feac3990",
899 => x"1a087a08",
900 => x"71317611",
901 => x"70565a57",
902 => x"5280d3f0",
903 => x"08519084",
904 => x"3fb00880",
905 => x"2effa738",
906 => x"b008901b",
907 => x"0cb00816",
908 => x"7a0c7794",
909 => x"1b0c7488",
910 => x"1b0c7456",
911 => x"fd993979",
912 => x"0858901a",
913 => x"08782783",
914 => x"38815475",
915 => x"75278438",
916 => x"73b33894",
917 => x"1a085675",
918 => x"752680d3",
919 => x"38755378",
920 => x"529c1a08",
921 => x"51a41a08",
922 => x"54732db0",
923 => x"0856b008",
924 => x"8024fd83",
925 => x"388c1a22",
926 => x"80c00754",
927 => x"738c1b23",
928 => x"ff54fed7",
929 => x"39755378",
930 => x"5277518d",
931 => x"d23f7908",
932 => x"167a0c79",
933 => x"5199a93f",
934 => x"b008802e",
935 => x"fcd9388c",
936 => x"1a2280c0",
937 => x"0754738c",
938 => x"1b23ff54",
939 => x"fead3974",
940 => x"75547953",
941 => x"7852568d",
942 => x"a63f881a",
943 => x"08753188",
944 => x"1b0c7908",
945 => x"157a0cfc",
946 => x"ae39f33d",
947 => x"0d7f618b",
948 => x"1170f806",
949 => x"5c55555e",
950 => x"72962683",
951 => x"38905980",
952 => x"7924747a",
953 => x"26075380",
954 => x"5472742e",
955 => x"09810680",
956 => x"cb387d51",
957 => x"8eac3f78",
958 => x"83f72680",
959 => x"c6387883",
960 => x"2a701010",
961 => x"1080dbac",
962 => x"058c1108",
963 => x"59595a76",
964 => x"782e83b0",
965 => x"38841708",
966 => x"fc06568c",
967 => x"17088818",
968 => x"08718c12",
969 => x"0c88120c",
970 => x"58751784",
971 => x"11088107",
972 => x"84120c53",
973 => x"7d518deb",
974 => x"3f881754",
975 => x"73b00c8f",
976 => x"3d0d0478",
977 => x"892a7983",
978 => x"2a5b5372",
979 => x"802ebf38",
980 => x"78862ab8",
981 => x"055a8473",
982 => x"27b43880",
983 => x"db135a94",
984 => x"7327ab38",
985 => x"788c2a80",
986 => x"ee055a80",
987 => x"d473279e",
988 => x"38788f2a",
989 => x"80f7055a",
990 => x"82d47327",
991 => x"91387892",
992 => x"2a80fc05",
993 => x"5a8ad473",
994 => x"27843880",
995 => x"fe5a7910",
996 => x"101080db",
997 => x"ac058c11",
998 => x"08585576",
999 => x"752ea338",
1000 => x"841708fc",
1001 => x"06707a31",
1002 => x"5556738f",
1003 => x"2488d538",
1004 => x"738025fe",
1005 => x"e6388c17",
1006 => x"08577675",
1007 => x"2e098106",
1008 => x"df38811a",
1009 => x"5a80dbbc",
1010 => x"08577680",
1011 => x"dbb42e82",
1012 => x"c0388417",
1013 => x"08fc0670",
1014 => x"7a315556",
1015 => x"738f2481",
1016 => x"f93880db",
1017 => x"b40b80db",
1018 => x"c00c80db",
1019 => x"b40b80db",
1020 => x"bc0c7380",
1021 => x"25feb238",
1022 => x"83ff7627",
1023 => x"83df3875",
1024 => x"892a7683",
1025 => x"2a555372",
1026 => x"802ebf38",
1027 => x"75862ab8",
1028 => x"05548473",
1029 => x"27b43880",
1030 => x"db135494",
1031 => x"7327ab38",
1032 => x"758c2a80",
1033 => x"ee055480",
1034 => x"d473279e",
1035 => x"38758f2a",
1036 => x"80f70554",
1037 => x"82d47327",
1038 => x"91387592",
1039 => x"2a80fc05",
1040 => x"548ad473",
1041 => x"27843880",
1042 => x"fe547310",
1043 => x"101080db",
1044 => x"ac058811",
1045 => x"08565874",
1046 => x"782e86cf",
1047 => x"38841508",
1048 => x"fc065375",
1049 => x"73278d38",
1050 => x"88150855",
1051 => x"74782e09",
1052 => x"8106ea38",
1053 => x"8c150880",
1054 => x"dbac0b84",
1055 => x"0508718c",
1056 => x"1a0c7688",
1057 => x"1a0c7888",
1058 => x"130c788c",
1059 => x"180c5d58",
1060 => x"7953807a",
1061 => x"2483e638",
1062 => x"72822c81",
1063 => x"712b5c53",
1064 => x"7a7c2681",
1065 => x"98387b7b",
1066 => x"06537282",
1067 => x"f13879fc",
1068 => x"0684055a",
1069 => x"7a10707d",
1070 => x"06545b72",
1071 => x"82e03884",
1072 => x"1a5af139",
1073 => x"88178c11",
1074 => x"08585876",
1075 => x"782e0981",
1076 => x"06fcc238",
1077 => x"821a5afd",
1078 => x"ec397817",
1079 => x"79810784",
1080 => x"190c7080",
1081 => x"dbc00c70",
1082 => x"80dbbc0c",
1083 => x"80dbb40b",
1084 => x"8c120c8c",
1085 => x"11088812",
1086 => x"0c748107",
1087 => x"84120c74",
1088 => x"1175710c",
1089 => x"51537d51",
1090 => x"8a993f88",
1091 => x"1754fcac",
1092 => x"3980dbac",
1093 => x"0b840508",
1094 => x"7a545c79",
1095 => x"8025fef8",
1096 => x"3882da39",
1097 => x"7a097c06",
1098 => x"7080dbac",
1099 => x"0b84050c",
1100 => x"5c7a105b",
1101 => x"7a7c2685",
1102 => x"387a85b8",
1103 => x"3880dbac",
1104 => x"0b880508",
1105 => x"70841208",
1106 => x"fc06707c",
1107 => x"317c7226",
1108 => x"8f722507",
1109 => x"57575c5d",
1110 => x"5572802e",
1111 => x"80db3879",
1112 => x"7a1680db",
1113 => x"a4081b90",
1114 => x"115a5557",
1115 => x"5b80dba0",
1116 => x"08ff2e88",
1117 => x"38a08f13",
1118 => x"e0800657",
1119 => x"76527d51",
1120 => x"91a73fb0",
1121 => x"0854b008",
1122 => x"ff2e9038",
1123 => x"b0087627",
1124 => x"82993874",
1125 => x"80dbac2e",
1126 => x"82913880",
1127 => x"dbac0b88",
1128 => x"05085584",
1129 => x"1508fc06",
1130 => x"707a317a",
1131 => x"72268f72",
1132 => x"25075255",
1133 => x"537283e6",
1134 => x"38747981",
1135 => x"0784170c",
1136 => x"79167080",
1137 => x"dbac0b88",
1138 => x"050c7581",
1139 => x"0784120c",
1140 => x"547e5257",
1141 => x"88cd3f88",
1142 => x"1754fae0",
1143 => x"3975832a",
1144 => x"70545480",
1145 => x"7424819b",
1146 => x"3872822c",
1147 => x"81712b80",
1148 => x"dbb00807",
1149 => x"7080dbac",
1150 => x"0b84050c",
1151 => x"75101010",
1152 => x"80dbac05",
1153 => x"88110858",
1154 => x"5a5d5377",
1155 => x"8c180c74",
1156 => x"88180c76",
1157 => x"88190c76",
1158 => x"8c160cfc",
1159 => x"f339797a",
1160 => x"10101080",
1161 => x"dbac0570",
1162 => x"57595d8c",
1163 => x"15085776",
1164 => x"752ea338",
1165 => x"841708fc",
1166 => x"06707a31",
1167 => x"5556738f",
1168 => x"2483ca38",
1169 => x"73802584",
1170 => x"81388c17",
1171 => x"08577675",
1172 => x"2e098106",
1173 => x"df388815",
1174 => x"811b7083",
1175 => x"06555b55",
1176 => x"72c9387c",
1177 => x"83065372",
1178 => x"802efdb8",
1179 => x"38ff1df8",
1180 => x"19595d88",
1181 => x"1808782e",
1182 => x"ea38fdb5",
1183 => x"39831a53",
1184 => x"fc963983",
1185 => x"1470822c",
1186 => x"81712b80",
1187 => x"dbb00807",
1188 => x"7080dbac",
1189 => x"0b84050c",
1190 => x"76101010",
1191 => x"80dbac05",
1192 => x"88110859",
1193 => x"5b5e5153",
1194 => x"fee13980",
1195 => x"daf00817",
1196 => x"58b00876",
1197 => x"2e818d38",
1198 => x"80dba008",
1199 => x"ff2e83ec",
1200 => x"38737631",
1201 => x"1880daf0",
1202 => x"0c738706",
1203 => x"70575372",
1204 => x"802e8838",
1205 => x"88733170",
1206 => x"15555676",
1207 => x"149fff06",
1208 => x"a0807131",
1209 => x"1770547f",
1210 => x"5357538e",
1211 => x"bc3fb008",
1212 => x"53b008ff",
1213 => x"2e81a038",
1214 => x"80daf008",
1215 => x"167080da",
1216 => x"f00c7475",
1217 => x"80dbac0b",
1218 => x"88050c74",
1219 => x"76311870",
1220 => x"81075155",
1221 => x"56587b80",
1222 => x"dbac2e83",
1223 => x"9c38798f",
1224 => x"2682cb38",
1225 => x"810b8415",
1226 => x"0c841508",
1227 => x"fc06707a",
1228 => x"317a7226",
1229 => x"8f722507",
1230 => x"52555372",
1231 => x"802efcf9",
1232 => x"3880db39",
1233 => x"b0089fff",
1234 => x"065372fe",
1235 => x"eb387780",
1236 => x"daf00c80",
1237 => x"dbac0b88",
1238 => x"05087b18",
1239 => x"81078412",
1240 => x"0c5580db",
1241 => x"9c087827",
1242 => x"86387780",
1243 => x"db9c0c80",
1244 => x"db980878",
1245 => x"27fcac38",
1246 => x"7780db98",
1247 => x"0c841508",
1248 => x"fc06707a",
1249 => x"317a7226",
1250 => x"8f722507",
1251 => x"52555372",
1252 => x"802efca5",
1253 => x"38883980",
1254 => x"745456fe",
1255 => x"db397d51",
1256 => x"85813f80",
1257 => x"0bb00c8f",
1258 => x"3d0d0473",
1259 => x"53807424",
1260 => x"a9387282",
1261 => x"2c81712b",
1262 => x"80dbb008",
1263 => x"077080db",
1264 => x"ac0b8405",
1265 => x"0c5d5377",
1266 => x"8c180c74",
1267 => x"88180c76",
1268 => x"88190c76",
1269 => x"8c160cf9",
1270 => x"b7398314",
1271 => x"70822c81",
1272 => x"712b80db",
1273 => x"b0080770",
1274 => x"80dbac0b",
1275 => x"84050c5e",
1276 => x"5153d439",
1277 => x"7b7b0653",
1278 => x"72fca338",
1279 => x"841a7b10",
1280 => x"5c5af139",
1281 => x"ff1a8111",
1282 => x"515af7b9",
1283 => x"39781779",
1284 => x"81078419",
1285 => x"0c8c1808",
1286 => x"88190871",
1287 => x"8c120c88",
1288 => x"120c5970",
1289 => x"80dbc00c",
1290 => x"7080dbbc",
1291 => x"0c80dbb4",
1292 => x"0b8c120c",
1293 => x"8c110888",
1294 => x"120c7481",
1295 => x"0784120c",
1296 => x"74117571",
1297 => x"0c5153f9",
1298 => x"bd397517",
1299 => x"84110881",
1300 => x"0784120c",
1301 => x"538c1708",
1302 => x"88180871",
1303 => x"8c120c88",
1304 => x"120c587d",
1305 => x"5183bc3f",
1306 => x"881754f5",
1307 => x"cf397284",
1308 => x"150cf41a",
1309 => x"f8067084",
1310 => x"1e088106",
1311 => x"07841e0c",
1312 => x"701d545b",
1313 => x"850b8414",
1314 => x"0c850b88",
1315 => x"140c8f7b",
1316 => x"27fdcf38",
1317 => x"881c527d",
1318 => x"5193ed3f",
1319 => x"80dbac0b",
1320 => x"88050880",
1321 => x"daf00859",
1322 => x"55fdb739",
1323 => x"7780daf0",
1324 => x"0c7380db",
1325 => x"a00cfc91",
1326 => x"39728415",
1327 => x"0cfda339",
1328 => x"fa3d0d7a",
1329 => x"79028805",
1330 => x"a7053356",
1331 => x"52538373",
1332 => x"278a3870",
1333 => x"83065271",
1334 => x"802ea838",
1335 => x"ff135372",
1336 => x"ff2e9738",
1337 => x"70335273",
1338 => x"722e9138",
1339 => x"8111ff14",
1340 => x"545172ff",
1341 => x"2e098106",
1342 => x"eb388051",
1343 => x"70b00c88",
1344 => x"3d0d0470",
1345 => x"72575583",
1346 => x"51758280",
1347 => x"2914ff12",
1348 => x"52567080",
1349 => x"25f33883",
1350 => x"7327bf38",
1351 => x"74087632",
1352 => x"7009f7fb",
1353 => x"fdff1206",
1354 => x"70f88482",
1355 => x"81800651",
1356 => x"51517080",
1357 => x"2e993874",
1358 => x"51805270",
1359 => x"33577377",
1360 => x"2effb938",
1361 => x"81118113",
1362 => x"53518372",
1363 => x"27ed38fc",
1364 => x"13841656",
1365 => x"53728326",
1366 => x"c3387451",
1367 => x"fefe39fa",
1368 => x"3d0d787a",
1369 => x"7c727272",
1370 => x"57575759",
1371 => x"56567476",
1372 => x"27b23876",
1373 => x"15517571",
1374 => x"27aa3870",
1375 => x"7717ff14",
1376 => x"54555371",
1377 => x"ff2e9638",
1378 => x"ff14ff14",
1379 => x"54547233",
1380 => x"7434ff12",
1381 => x"5271ff2e",
1382 => x"098106ec",
1383 => x"3875b00c",
1384 => x"883d0d04",
1385 => x"768f2697",
1386 => x"38ff1252",
1387 => x"71ff2eed",
1388 => x"38727081",
1389 => x"05543374",
1390 => x"70810556",
1391 => x"34eb3974",
1392 => x"76078306",
1393 => x"5170e238",
1394 => x"75755451",
1395 => x"72708405",
1396 => x"54087170",
1397 => x"8405530c",
1398 => x"72708405",
1399 => x"54087170",
1400 => x"8405530c",
1401 => x"72708405",
1402 => x"54087170",
1403 => x"8405530c",
1404 => x"72708405",
1405 => x"54087170",
1406 => x"8405530c",
1407 => x"f0125271",
1408 => x"8f26c938",
1409 => x"83722795",
1410 => x"38727084",
1411 => x"05540871",
1412 => x"70840553",
1413 => x"0cfc1252",
1414 => x"718326ed",
1415 => x"387054ff",
1416 => x"88390404",
1417 => x"ef3d0d63",
1418 => x"6567405d",
1419 => x"427b802e",
1420 => x"84f93861",
1421 => x"51ec3ff8",
1422 => x"1c708412",
1423 => x"0870fc06",
1424 => x"70628b05",
1425 => x"70f80641",
1426 => x"59455b5c",
1427 => x"41579674",
1428 => x"2782c338",
1429 => x"807b247e",
1430 => x"7c260759",
1431 => x"80547874",
1432 => x"2e098106",
1433 => x"82a93877",
1434 => x"7b2581fc",
1435 => x"38771780",
1436 => x"dbac0b88",
1437 => x"05085e56",
1438 => x"7c762e84",
1439 => x"bd388416",
1440 => x"0870fe06",
1441 => x"17841108",
1442 => x"81065155",
1443 => x"5573828b",
1444 => x"3874fc06",
1445 => x"597c762e",
1446 => x"84dd3877",
1447 => x"195f7e7b",
1448 => x"2581fd38",
1449 => x"79810654",
1450 => x"7382bf38",
1451 => x"76770831",
1452 => x"841108fc",
1453 => x"06565a75",
1454 => x"802e9138",
1455 => x"7c762e84",
1456 => x"ea387419",
1457 => x"1859787b",
1458 => x"25848938",
1459 => x"79802e82",
1460 => x"99387715",
1461 => x"567a7624",
1462 => x"8290388c",
1463 => x"1a08881b",
1464 => x"08718c12",
1465 => x"0c88120c",
1466 => x"55797659",
1467 => x"57881761",
1468 => x"fc055759",
1469 => x"75a42685",
1470 => x"ef387b79",
1471 => x"55559376",
1472 => x"2780c938",
1473 => x"7b708405",
1474 => x"5d087c56",
1475 => x"790c7470",
1476 => x"84055608",
1477 => x"8c180c90",
1478 => x"17549b76",
1479 => x"27ae3874",
1480 => x"70840556",
1481 => x"08740c74",
1482 => x"70840556",
1483 => x"0894180c",
1484 => x"981754a3",
1485 => x"76279538",
1486 => x"74708405",
1487 => x"5608740c",
1488 => x"74708405",
1489 => x"56089c18",
1490 => x"0ca01754",
1491 => x"74708405",
1492 => x"56087470",
1493 => x"8405560c",
1494 => x"74708405",
1495 => x"56087470",
1496 => x"8405560c",
1497 => x"7408740c",
1498 => x"777b3156",
1499 => x"758f2680",
1500 => x"c9388417",
1501 => x"08810678",
1502 => x"0784180c",
1503 => x"77178411",
1504 => x"08810784",
1505 => x"120c5461",
1506 => x"51fd983f",
1507 => x"88175473",
1508 => x"b00c933d",
1509 => x"0d04905b",
1510 => x"fdba3978",
1511 => x"56fe8539",
1512 => x"8c160888",
1513 => x"1708718c",
1514 => x"120c8812",
1515 => x"0c557e70",
1516 => x"7c315758",
1517 => x"8f7627ff",
1518 => x"b9387a17",
1519 => x"84180881",
1520 => x"067c0784",
1521 => x"190c7681",
1522 => x"0784120c",
1523 => x"76118411",
1524 => x"08810784",
1525 => x"120c5588",
1526 => x"05526151",
1527 => x"8daa3f61",
1528 => x"51fcc03f",
1529 => x"881754ff",
1530 => x"a6397d52",
1531 => x"6151edda",
1532 => x"3fb00859",
1533 => x"b008802e",
1534 => x"81a338b0",
1535 => x"08f80560",
1536 => x"840508fe",
1537 => x"06610555",
1538 => x"5776742e",
1539 => x"83e638fc",
1540 => x"185675a4",
1541 => x"2681aa38",
1542 => x"7bb00855",
1543 => x"55937627",
1544 => x"80d83874",
1545 => x"70840556",
1546 => x"08b00870",
1547 => x"8405b00c",
1548 => x"0cb00875",
1549 => x"70840557",
1550 => x"08717084",
1551 => x"05530c54",
1552 => x"9b7627b6",
1553 => x"38747084",
1554 => x"05560874",
1555 => x"70840556",
1556 => x"0c747084",
1557 => x"05560874",
1558 => x"70840556",
1559 => x"0ca37627",
1560 => x"99387470",
1561 => x"84055608",
1562 => x"74708405",
1563 => x"560c7470",
1564 => x"84055608",
1565 => x"74708405",
1566 => x"560c7470",
1567 => x"84055608",
1568 => x"74708405",
1569 => x"560c7470",
1570 => x"84055608",
1571 => x"74708405",
1572 => x"560c7408",
1573 => x"740c7b52",
1574 => x"61518bec",
1575 => x"3f6151fb",
1576 => x"823f7854",
1577 => x"73b00c93",
1578 => x"3d0d047d",
1579 => x"526151ec",
1580 => x"993fb008",
1581 => x"b00c933d",
1582 => x"0d048416",
1583 => x"0855fbd1",
1584 => x"3975537b",
1585 => x"52b00851",
1586 => x"dfdc3f7b",
1587 => x"5261518b",
1588 => x"b73fca39",
1589 => x"8c160888",
1590 => x"1708718c",
1591 => x"120c8812",
1592 => x"0c558c1a",
1593 => x"08881b08",
1594 => x"718c120c",
1595 => x"88120c55",
1596 => x"79795957",
1597 => x"fbf73977",
1598 => x"19901c55",
1599 => x"55737524",
1600 => x"fba2387a",
1601 => x"177080db",
1602 => x"ac0b8805",
1603 => x"0c757c31",
1604 => x"81078412",
1605 => x"0c5d8417",
1606 => x"0881067b",
1607 => x"0784180c",
1608 => x"6151f9ff",
1609 => x"3f881754",
1610 => x"fce53974",
1611 => x"1918901c",
1612 => x"555d737d",
1613 => x"24fb9538",
1614 => x"8c1a0888",
1615 => x"1b08718c",
1616 => x"120c8812",
1617 => x"0c55881a",
1618 => x"61fc0557",
1619 => x"5975a426",
1620 => x"81ae387b",
1621 => x"79555593",
1622 => x"762780c9",
1623 => x"387b7084",
1624 => x"055d087c",
1625 => x"56790c74",
1626 => x"70840556",
1627 => x"088c1b0c",
1628 => x"901a549b",
1629 => x"7627ae38",
1630 => x"74708405",
1631 => x"5608740c",
1632 => x"74708405",
1633 => x"5608941b",
1634 => x"0c981a54",
1635 => x"a3762795",
1636 => x"38747084",
1637 => x"05560874",
1638 => x"0c747084",
1639 => x"0556089c",
1640 => x"1b0ca01a",
1641 => x"54747084",
1642 => x"05560874",
1643 => x"70840556",
1644 => x"0c747084",
1645 => x"05560874",
1646 => x"70840556",
1647 => x"0c740874",
1648 => x"0c7a1a70",
1649 => x"80dbac0b",
1650 => x"88050c7d",
1651 => x"7c318107",
1652 => x"84120c54",
1653 => x"841a0881",
1654 => x"067b0784",
1655 => x"1b0c6151",
1656 => x"f8c13f78",
1657 => x"54fdbd39",
1658 => x"75537b52",
1659 => x"7851ddb6",
1660 => x"3ffaf539",
1661 => x"841708fc",
1662 => x"06186058",
1663 => x"58fae939",
1664 => x"75537b52",
1665 => x"7851dd9e",
1666 => x"3f7a1a70",
1667 => x"80dbac0b",
1668 => x"88050c7d",
1669 => x"7c318107",
1670 => x"84120c54",
1671 => x"841a0881",
1672 => x"067b0784",
1673 => x"1b0cffb6",
1674 => x"39fd3d0d",
1675 => x"800b80e3",
1676 => x"e40c7651",
1677 => x"96d33fb0",
1678 => x"0853b008",
1679 => x"ff2e8838",
1680 => x"72b00c85",
1681 => x"3d0d0480",
1682 => x"e3e40854",
1683 => x"73802ef0",
1684 => x"38757471",
1685 => x"0c5272b0",
1686 => x"0c853d0d",
1687 => x"04fa3d0d",
1688 => x"7880d3f0",
1689 => x"085455b8",
1690 => x"1308802e",
1691 => x"81b5388c",
1692 => x"15227083",
1693 => x"ffff0670",
1694 => x"832a8132",
1695 => x"70810651",
1696 => x"55555672",
1697 => x"802e80dc",
1698 => x"3873842a",
1699 => x"81328106",
1700 => x"57ff5376",
1701 => x"80f63873",
1702 => x"822a7081",
1703 => x"06515372",
1704 => x"802eb938",
1705 => x"b0150854",
1706 => x"73802e9c",
1707 => x"3880c015",
1708 => x"5373732e",
1709 => x"8f387352",
1710 => x"80d3f008",
1711 => x"5187c93f",
1712 => x"8c152256",
1713 => x"76b0160c",
1714 => x"75db0653",
1715 => x"728c1623",
1716 => x"800b8416",
1717 => x"0c901508",
1718 => x"750c7256",
1719 => x"75880753",
1720 => x"728c1623",
1721 => x"90150880",
1722 => x"2e80c038",
1723 => x"8c152270",
1724 => x"81065553",
1725 => x"739d3872",
1726 => x"812a7081",
1727 => x"06515372",
1728 => x"85389415",
1729 => x"08547388",
1730 => x"160c8053",
1731 => x"72b00c88",
1732 => x"3d0d0480",
1733 => x"0b88160c",
1734 => x"94150830",
1735 => x"98160c80",
1736 => x"53ea3972",
1737 => x"5182fb3f",
1738 => x"fec53974",
1739 => x"518ce83f",
1740 => x"8c152270",
1741 => x"81065553",
1742 => x"73802eff",
1743 => x"ba38d439",
1744 => x"f83d0d7a",
1745 => x"5877802e",
1746 => x"81993880",
1747 => x"d3f00854",
1748 => x"b8140880",
1749 => x"2e80ed38",
1750 => x"8c182270",
1751 => x"902b7090",
1752 => x"2c70832a",
1753 => x"81328106",
1754 => x"5c515754",
1755 => x"7880cd38",
1756 => x"90180857",
1757 => x"76802e80",
1758 => x"c3387708",
1759 => x"77317779",
1760 => x"0c768306",
1761 => x"7a585555",
1762 => x"73853894",
1763 => x"18085675",
1764 => x"88190c80",
1765 => x"7525a538",
1766 => x"74537652",
1767 => x"9c180851",
1768 => x"a4180854",
1769 => x"732d800b",
1770 => x"b0082580",
1771 => x"c938b008",
1772 => x"1775b008",
1773 => x"31565774",
1774 => x"8024dd38",
1775 => x"800bb00c",
1776 => x"8a3d0d04",
1777 => x"735181da",
1778 => x"3f8c1822",
1779 => x"70902b70",
1780 => x"902c7083",
1781 => x"2a813281",
1782 => x"065c5157",
1783 => x"5478dd38",
1784 => x"ff8e39b6",
1785 => x"c05280d3",
1786 => x"f0085189",
1787 => x"f13fb008",
1788 => x"b00c8a3d",
1789 => x"0d048c18",
1790 => x"2280c007",
1791 => x"54738c19",
1792 => x"23ff0bb0",
1793 => x"0c8a3d0d",
1794 => x"04803d0d",
1795 => x"72518071",
1796 => x"0c800b84",
1797 => x"120c800b",
1798 => x"88120c02",
1799 => x"8e05228c",
1800 => x"12230292",
1801 => x"05228e12",
1802 => x"23800b90",
1803 => x"120c800b",
1804 => x"94120c80",
1805 => x"0b98120c",
1806 => x"709c120c",
1807 => x"80c6a80b",
1808 => x"a0120c80",
1809 => x"c6f40ba4",
1810 => x"120c80c7",
1811 => x"f00ba812",
1812 => x"0c80c8c1",
1813 => x"0bac120c",
1814 => x"823d0d04",
1815 => x"fa3d0d79",
1816 => x"7080dc29",
1817 => x"8c11547a",
1818 => x"535657e4",
1819 => x"dd3fb008",
1820 => x"b0085556",
1821 => x"b008802e",
1822 => x"a238b008",
1823 => x"8c055480",
1824 => x"0bb0080c",
1825 => x"76b00884",
1826 => x"050c73b0",
1827 => x"0888050c",
1828 => x"74538052",
1829 => x"73518c81",
1830 => x"3f755473",
1831 => x"b00c883d",
1832 => x"0d04fc3d",
1833 => x"0d76bbb5",
1834 => x"0bbc120c",
1835 => x"55810bb8",
1836 => x"160c800b",
1837 => x"84dc160c",
1838 => x"830b84e0",
1839 => x"160c84e8",
1840 => x"1584e416",
1841 => x"0c745480",
1842 => x"53845284",
1843 => x"150851fe",
1844 => x"b83f7454",
1845 => x"81538952",
1846 => x"88150851",
1847 => x"feab3f74",
1848 => x"5482538a",
1849 => x"528c1508",
1850 => x"51fe9e3f",
1851 => x"863d0d04",
1852 => x"f93d0d79",
1853 => x"80d3f008",
1854 => x"5457b813",
1855 => x"08802e80",
1856 => x"c83884dc",
1857 => x"13568816",
1858 => x"08841708",
1859 => x"ff055555",
1860 => x"8074249f",
1861 => x"388c1522",
1862 => x"70902b70",
1863 => x"902c5154",
1864 => x"5872802e",
1865 => x"80ca3880",
1866 => x"dc15ff15",
1867 => x"55557380",
1868 => x"25e33875",
1869 => x"08537280",
1870 => x"2e9f3872",
1871 => x"56881608",
1872 => x"841708ff",
1873 => x"055555c8",
1874 => x"397251fe",
1875 => x"d53f80d3",
1876 => x"f00884dc",
1877 => x"0556ffae",
1878 => x"39845276",
1879 => x"51fdfd3f",
1880 => x"b008760c",
1881 => x"b008802e",
1882 => x"80c038b0",
1883 => x"0856ce39",
1884 => x"810b8c16",
1885 => x"2372750c",
1886 => x"7288160c",
1887 => x"7284160c",
1888 => x"7290160c",
1889 => x"7294160c",
1890 => x"7298160c",
1891 => x"ff0b8e16",
1892 => x"2372b016",
1893 => x"0c72b416",
1894 => x"0c7280c4",
1895 => x"160c7280",
1896 => x"c8160c74",
1897 => x"b00c893d",
1898 => x"0d048c77",
1899 => x"0c800bb0",
1900 => x"0c893d0d",
1901 => x"04ff3d0d",
1902 => x"b6c05273",
1903 => x"51869f3f",
1904 => x"833d0d04",
1905 => x"803d0d80",
1906 => x"d3f00851",
1907 => x"e83f823d",
1908 => x"0d04fb3d",
1909 => x"0d777052",
1910 => x"56f0c73f",
1911 => x"80dbac0b",
1912 => x"88050884",
1913 => x"1108fc06",
1914 => x"707b319f",
1915 => x"ef05e080",
1916 => x"06e08005",
1917 => x"565653a0",
1918 => x"80742494",
1919 => x"38805275",
1920 => x"51f8a63f",
1921 => x"80dbb408",
1922 => x"155372b0",
1923 => x"082e8f38",
1924 => x"7551f08f",
1925 => x"3f805372",
1926 => x"b00c873d",
1927 => x"0d047330",
1928 => x"527551f8",
1929 => x"843fb008",
1930 => x"ff2ea838",
1931 => x"80dbac0b",
1932 => x"88050875",
1933 => x"75318107",
1934 => x"84120c53",
1935 => x"80daf008",
1936 => x"743180da",
1937 => x"f00c7551",
1938 => x"efd93f81",
1939 => x"0bb00c87",
1940 => x"3d0d0480",
1941 => x"527551f7",
1942 => x"d03f80db",
1943 => x"ac0b8805",
1944 => x"08b00871",
1945 => x"3156538f",
1946 => x"7525ffa4",
1947 => x"38b00880",
1948 => x"dba00831",
1949 => x"80daf00c",
1950 => x"74810784",
1951 => x"140c7551",
1952 => x"efa13f80",
1953 => x"53ff9039",
1954 => x"f63d0d7c",
1955 => x"7e545b72",
1956 => x"802e8283",
1957 => x"387a51ef",
1958 => x"893ff813",
1959 => x"84110870",
1960 => x"fe067013",
1961 => x"841108fc",
1962 => x"065d5859",
1963 => x"545880db",
1964 => x"b408752e",
1965 => x"82de3878",
1966 => x"84160c80",
1967 => x"73810654",
1968 => x"5a727a2e",
1969 => x"81d53878",
1970 => x"15841108",
1971 => x"81065153",
1972 => x"72a03878",
1973 => x"17577981",
1974 => x"e6388815",
1975 => x"08537280",
1976 => x"dbb42e82",
1977 => x"f9388c15",
1978 => x"08708c15",
1979 => x"0c738812",
1980 => x"0c567681",
1981 => x"0784190c",
1982 => x"76187771",
1983 => x"0c537981",
1984 => x"913883ff",
1985 => x"772781c8",
1986 => x"3876892a",
1987 => x"77832a56",
1988 => x"5372802e",
1989 => x"bf387686",
1990 => x"2ab80555",
1991 => x"847327b4",
1992 => x"3880db13",
1993 => x"55947327",
1994 => x"ab38768c",
1995 => x"2a80ee05",
1996 => x"5580d473",
1997 => x"279e3876",
1998 => x"8f2a80f7",
1999 => x"055582d4",
2000 => x"73279138",
2001 => x"76922a80",
2002 => x"fc05558a",
2003 => x"d4732784",
2004 => x"3880fe55",
2005 => x"74101010",
2006 => x"80dbac05",
2007 => x"88110855",
2008 => x"5673762e",
2009 => x"82b33884",
2010 => x"1408fc06",
2011 => x"53767327",
2012 => x"8d388814",
2013 => x"08547376",
2014 => x"2e098106",
2015 => x"ea388c14",
2016 => x"08708c1a",
2017 => x"0c74881a",
2018 => x"0c788812",
2019 => x"0c56778c",
2020 => x"150c7a51",
2021 => x"ed8d3f8c",
2022 => x"3d0d0477",
2023 => x"08787131",
2024 => x"59770588",
2025 => x"19085457",
2026 => x"7280dbb4",
2027 => x"2e80e038",
2028 => x"8c180870",
2029 => x"8c150c73",
2030 => x"88120c56",
2031 => x"fe893988",
2032 => x"15088c16",
2033 => x"08708c13",
2034 => x"0c578817",
2035 => x"0cfea339",
2036 => x"76832a70",
2037 => x"54558075",
2038 => x"24819838",
2039 => x"72822c81",
2040 => x"712b80db",
2041 => x"b0080780",
2042 => x"dbac0b84",
2043 => x"050c5374",
2044 => x"10101080",
2045 => x"dbac0588",
2046 => x"11085556",
2047 => x"758c190c",
2048 => x"7388190c",
2049 => x"7788170c",
2050 => x"778c150c",
2051 => x"ff843981",
2052 => x"5afdb439",
2053 => x"78177381",
2054 => x"06545772",
2055 => x"98387708",
2056 => x"78713159",
2057 => x"77058c19",
2058 => x"08881a08",
2059 => x"718c120c",
2060 => x"88120c57",
2061 => x"57768107",
2062 => x"84190c77",
2063 => x"80dbac0b",
2064 => x"88050c80",
2065 => x"dba80877",
2066 => x"26fec738",
2067 => x"80dba408",
2068 => x"527a51fa",
2069 => x"fd3f7a51",
2070 => x"ebc93ffe",
2071 => x"ba398178",
2072 => x"8c150c78",
2073 => x"88150c73",
2074 => x"8c1a0c73",
2075 => x"881a0c5a",
2076 => x"fd803983",
2077 => x"1570822c",
2078 => x"81712b80",
2079 => x"dbb00807",
2080 => x"80dbac0b",
2081 => x"84050c51",
2082 => x"53741010",
2083 => x"1080dbac",
2084 => x"05881108",
2085 => x"5556fee4",
2086 => x"39745380",
2087 => x"7524a738",
2088 => x"72822c81",
2089 => x"712b80db",
2090 => x"b0080780",
2091 => x"dbac0b84",
2092 => x"050c5375",
2093 => x"8c190c73",
2094 => x"88190c77",
2095 => x"88170c77",
2096 => x"8c150cfd",
2097 => x"cd398315",
2098 => x"70822c81",
2099 => x"712b80db",
2100 => x"b0080780",
2101 => x"dbac0b84",
2102 => x"050c5153",
2103 => x"d639f93d",
2104 => x"0d797b58",
2105 => x"53800b80",
2106 => x"d3f00853",
2107 => x"5672722e",
2108 => x"80c03884",
2109 => x"dc135574",
2110 => x"762eb738",
2111 => x"88150884",
2112 => x"1608ff05",
2113 => x"54548073",
2114 => x"249d388c",
2115 => x"14227090",
2116 => x"2b70902c",
2117 => x"51535871",
2118 => x"80d83880",
2119 => x"dc14ff14",
2120 => x"54547280",
2121 => x"25e53874",
2122 => x"085574d0",
2123 => x"3880d3f0",
2124 => x"085284dc",
2125 => x"12557480",
2126 => x"2eb13888",
2127 => x"15088416",
2128 => x"08ff0554",
2129 => x"54807324",
2130 => x"9c388c14",
2131 => x"2270902b",
2132 => x"70902c51",
2133 => x"535871ad",
2134 => x"3880dc14",
2135 => x"ff145454",
2136 => x"728025e6",
2137 => x"38740855",
2138 => x"74d13875",
2139 => x"b00c893d",
2140 => x"0d047351",
2141 => x"762d75b0",
2142 => x"080780dc",
2143 => x"15ff1555",
2144 => x"5556ff9e",
2145 => x"39735176",
2146 => x"2d75b008",
2147 => x"0780dc15",
2148 => x"ff155555",
2149 => x"56ca39ea",
2150 => x"3d0d688c",
2151 => x"11227081",
2152 => x"2a810657",
2153 => x"58567480",
2154 => x"e4388e16",
2155 => x"2270902b",
2156 => x"70902c51",
2157 => x"55588074",
2158 => x"24b13898",
2159 => x"3dc40553",
2160 => x"735280d3",
2161 => x"f0085186",
2162 => x"803f800b",
2163 => x"b0082497",
2164 => x"387983e0",
2165 => x"80065473",
2166 => x"80c0802e",
2167 => x"818f3873",
2168 => x"8280802e",
2169 => x"8191388c",
2170 => x"16225776",
2171 => x"90800754",
2172 => x"738c1723",
2173 => x"88805280",
2174 => x"d3f00851",
2175 => x"d9cc3fb0",
2176 => x"089d388c",
2177 => x"16228207",
2178 => x"54738c17",
2179 => x"2380c316",
2180 => x"70770c90",
2181 => x"170c810b",
2182 => x"94170c98",
2183 => x"3d0d0480",
2184 => x"d3f008bb",
2185 => x"b50bbc12",
2186 => x"0c548c16",
2187 => x"22818007",
2188 => x"54738c17",
2189 => x"23b00876",
2190 => x"0cb00890",
2191 => x"170c8880",
2192 => x"0b94170c",
2193 => x"74802ed3",
2194 => x"388e1622",
2195 => x"70902b70",
2196 => x"902c5355",
2197 => x"588ca13f",
2198 => x"b008802e",
2199 => x"ffbd388c",
2200 => x"16228107",
2201 => x"54738c17",
2202 => x"23983d0d",
2203 => x"04810b8c",
2204 => x"17225855",
2205 => x"fef539a8",
2206 => x"160880c7",
2207 => x"f02e0981",
2208 => x"06fee438",
2209 => x"8c162288",
2210 => x"80075473",
2211 => x"8c172388",
2212 => x"800b80cc",
2213 => x"170cfedc",
2214 => x"39fc3d0d",
2215 => x"76797102",
2216 => x"8c059f05",
2217 => x"33575553",
2218 => x"55837227",
2219 => x"8a387483",
2220 => x"06517080",
2221 => x"2ea238ff",
2222 => x"125271ff",
2223 => x"2e933873",
2224 => x"73708105",
2225 => x"5534ff12",
2226 => x"5271ff2e",
2227 => x"098106ef",
2228 => x"3874b00c",
2229 => x"863d0d04",
2230 => x"7474882b",
2231 => x"75077071",
2232 => x"902b0751",
2233 => x"54518f72",
2234 => x"27a53872",
2235 => x"71708405",
2236 => x"530c7271",
2237 => x"70840553",
2238 => x"0c727170",
2239 => x"8405530c",
2240 => x"72717084",
2241 => x"05530cf0",
2242 => x"1252718f",
2243 => x"26dd3883",
2244 => x"72279038",
2245 => x"72717084",
2246 => x"05530cfc",
2247 => x"12527183",
2248 => x"26f23870",
2249 => x"53ff9039",
2250 => x"f93d0d79",
2251 => x"7c557b54",
2252 => x"8e112270",
2253 => x"902b7090",
2254 => x"2c555780",
2255 => x"d3f00853",
2256 => x"585683f3",
2257 => x"3fb00857",
2258 => x"800bb008",
2259 => x"24933880",
2260 => x"d01608b0",
2261 => x"080580d0",
2262 => x"170c76b0",
2263 => x"0c893d0d",
2264 => x"048c1622",
2265 => x"83dfff06",
2266 => x"55748c17",
2267 => x"2376b00c",
2268 => x"893d0d04",
2269 => x"fa3d0d78",
2270 => x"8c112270",
2271 => x"882a7081",
2272 => x"06515758",
2273 => x"5674a938",
2274 => x"8c162283",
2275 => x"dfff0655",
2276 => x"748c1723",
2277 => x"7a547953",
2278 => x"8e162270",
2279 => x"902b7090",
2280 => x"2c545680",
2281 => x"d3f00852",
2282 => x"5681b23f",
2283 => x"883d0d04",
2284 => x"82548053",
2285 => x"8e162270",
2286 => x"902b7090",
2287 => x"2c545680",
2288 => x"d3f00852",
2289 => x"5782b83f",
2290 => x"8c162283",
2291 => x"dfff0655",
2292 => x"748c1723",
2293 => x"7a547953",
2294 => x"8e162270",
2295 => x"902b7090",
2296 => x"2c545680",
2297 => x"d3f00852",
2298 => x"5680f23f",
2299 => x"883d0d04",
2300 => x"f93d0d79",
2301 => x"7c557b54",
2302 => x"8e112270",
2303 => x"902b7090",
2304 => x"2c555780",
2305 => x"d3f00853",
2306 => x"585681f3",
2307 => x"3fb00857",
2308 => x"b008ff2e",
2309 => x"99388c16",
2310 => x"22a08007",
2311 => x"55748c17",
2312 => x"23b00880",
2313 => x"d0170c76",
2314 => x"b00c893d",
2315 => x"0d048c16",
2316 => x"2283dfff",
2317 => x"0655748c",
2318 => x"172376b0",
2319 => x"0c893d0d",
2320 => x"04fe3d0d",
2321 => x"748e1122",
2322 => x"70902b70",
2323 => x"902c5551",
2324 => x"515380d3",
2325 => x"f00851bd",
2326 => x"3f843d0d",
2327 => x"04fb3d0d",
2328 => x"800b80e3",
2329 => x"e40c7a53",
2330 => x"79527851",
2331 => x"839a3fb0",
2332 => x"0855b008",
2333 => x"ff2e8838",
2334 => x"74b00c87",
2335 => x"3d0d0480",
2336 => x"e3e40856",
2337 => x"75802ef0",
2338 => x"38777671",
2339 => x"0c5474b0",
2340 => x"0c873d0d",
2341 => x"04fd3d0d",
2342 => x"800b80e3",
2343 => x"e40c7651",
2344 => x"84ef3fb0",
2345 => x"0853b008",
2346 => x"ff2e8838",
2347 => x"72b00c85",
2348 => x"3d0d0480",
2349 => x"e3e40854",
2350 => x"73802ef0",
2351 => x"38757471",
2352 => x"0c5272b0",
2353 => x"0c853d0d",
2354 => x"04fc3d0d",
2355 => x"800b80e3",
2356 => x"e40c7852",
2357 => x"775186d7",
2358 => x"3fb00854",
2359 => x"b008ff2e",
2360 => x"883873b0",
2361 => x"0c863d0d",
2362 => x"0480e3e4",
2363 => x"08557480",
2364 => x"2ef03876",
2365 => x"75710c53",
2366 => x"73b00c86",
2367 => x"3d0d04fb",
2368 => x"3d0d800b",
2369 => x"80e3e40c",
2370 => x"7a537952",
2371 => x"785184b3",
2372 => x"3fb00855",
2373 => x"b008ff2e",
2374 => x"883874b0",
2375 => x"0c873d0d",
2376 => x"0480e3e4",
2377 => x"08567580",
2378 => x"2ef03877",
2379 => x"76710c54",
2380 => x"74b00c87",
2381 => x"3d0d04fb",
2382 => x"3d0d800b",
2383 => x"80e3e40c",
2384 => x"7a537952",
2385 => x"785182b8",
2386 => x"3fb00855",
2387 => x"b008ff2e",
2388 => x"883874b0",
2389 => x"0c873d0d",
2390 => x"0480e3e4",
2391 => x"08567580",
2392 => x"2ef03877",
2393 => x"76710c54",
2394 => x"74b00c87",
2395 => x"3d0d0481",
2396 => x"0bb00c04",
2397 => x"803d0d72",
2398 => x"812e8938",
2399 => x"800bb00c",
2400 => x"823d0d04",
2401 => x"735180fa",
2402 => x"3ffe3d0d",
2403 => x"80e3dc08",
2404 => x"51708a38",
2405 => x"80e3e870",
2406 => x"80e3dc0c",
2407 => x"51707512",
2408 => x"5252ff53",
2409 => x"7087fb80",
2410 => x"80268838",
2411 => x"7080e3dc",
2412 => x"0c715372",
2413 => x"b00c843d",
2414 => x"0d04fd3d",
2415 => x"0d800b80",
2416 => x"d3e40854",
2417 => x"5472812e",
2418 => x"9d387380",
2419 => x"e3e00cff",
2420 => x"be953fff",
2421 => x"bcaa3f80",
2422 => x"e3b45281",
2423 => x"51c0bd3f",
2424 => x"b0085185",
2425 => x"ca3f7280",
2426 => x"e3e00cff",
2427 => x"bdf93fff",
2428 => x"bc8e3f80",
2429 => x"e3b45281",
2430 => x"51c0a13f",
2431 => x"b0085185",
2432 => x"ae3f00ff",
2433 => x"3900ff39",
2434 => x"f53d0d7e",
2435 => x"6080e3e0",
2436 => x"08705b58",
2437 => x"5b5b7580",
2438 => x"c538777a",
2439 => x"25a23877",
2440 => x"1b703370",
2441 => x"81ff0658",
2442 => x"5859758a",
2443 => x"2e993876",
2444 => x"81ff0651",
2445 => x"ffbd8f3f",
2446 => x"81185879",
2447 => x"7824e038",
2448 => x"79b00c8d",
2449 => x"3d0d048d",
2450 => x"51ffbcfa",
2451 => x"3f783370",
2452 => x"81ff0652",
2453 => x"57ffbcee",
2454 => x"3f811858",
2455 => x"de397955",
2456 => x"7a547d53",
2457 => x"85528d3d",
2458 => x"fc0551ff",
2459 => x"bbd43fb0",
2460 => x"085684b4",
2461 => x"3f7bb008",
2462 => x"0c75b00c",
2463 => x"8d3d0d04",
2464 => x"f63d0d7d",
2465 => x"7f80e3e0",
2466 => x"08705b58",
2467 => x"5a5a7580",
2468 => x"c4387779",
2469 => x"25b638ff",
2470 => x"bc873fb0",
2471 => x"0881ff06",
2472 => x"708d3270",
2473 => x"30709f2a",
2474 => x"51515757",
2475 => x"768a2e80",
2476 => x"c6387580",
2477 => x"2e80c038",
2478 => x"771a5676",
2479 => x"76347651",
2480 => x"ffbc833f",
2481 => x"81185878",
2482 => x"7824cc38",
2483 => x"775675b0",
2484 => x"0c8c3d0d",
2485 => x"04785579",
2486 => x"547c5384",
2487 => x"528c3dfc",
2488 => x"0551ffba",
2489 => x"dd3fb008",
2490 => x"5683bd3f",
2491 => x"7ab0080c",
2492 => x"75b00c8c",
2493 => x"3d0d0477",
2494 => x"1a568a76",
2495 => x"34811858",
2496 => x"8d51ffbb",
2497 => x"c13f8a51",
2498 => x"ffbbbb3f",
2499 => x"7756ffbe",
2500 => x"39fb3d0d",
2501 => x"80e3e008",
2502 => x"70565473",
2503 => x"883874b0",
2504 => x"0c873d0d",
2505 => x"04775383",
2506 => x"52873dfc",
2507 => x"0551ffba",
2508 => x"913fb008",
2509 => x"5482f13f",
2510 => x"75b0080c",
2511 => x"73b00c87",
2512 => x"3d0d04fa",
2513 => x"3d0d80e3",
2514 => x"e008802e",
2515 => x"a3387a55",
2516 => x"79547853",
2517 => x"8652883d",
2518 => x"fc0551ff",
2519 => x"b9e43fb0",
2520 => x"085682c4",
2521 => x"3f76b008",
2522 => x"0c75b00c",
2523 => x"883d0d04",
2524 => x"82b63f9d",
2525 => x"0bb0080c",
2526 => x"ff0bb00c",
2527 => x"883d0d04",
2528 => x"fb3d0d77",
2529 => x"79565680",
2530 => x"70545473",
2531 => x"75259f38",
2532 => x"74101010",
2533 => x"f8055272",
2534 => x"16703370",
2535 => x"742b7607",
2536 => x"8116f816",
2537 => x"56565651",
2538 => x"51747324",
2539 => x"ea3873b0",
2540 => x"0c873d0d",
2541 => x"04fc3d0d",
2542 => x"76785555",
2543 => x"bc538052",
2544 => x"7351f5d5",
2545 => x"3f845274",
2546 => x"51ffb53f",
2547 => x"b0087423",
2548 => x"84528415",
2549 => x"51ffa93f",
2550 => x"b0088215",
2551 => x"23845288",
2552 => x"1551ff9c",
2553 => x"3fb00884",
2554 => x"150c8452",
2555 => x"8c1551ff",
2556 => x"8f3fb008",
2557 => x"88152384",
2558 => x"52901551",
2559 => x"ff823fb0",
2560 => x"088a1523",
2561 => x"84529415",
2562 => x"51fef53f",
2563 => x"b0088c15",
2564 => x"23845298",
2565 => x"1551fee8",
2566 => x"3fb0088e",
2567 => x"15238852",
2568 => x"9c1551fe",
2569 => x"db3fb008",
2570 => x"90150c86",
2571 => x"3d0d04e9",
2572 => x"3d0d6a80",
2573 => x"e3e00857",
2574 => x"57759338",
2575 => x"80c0800b",
2576 => x"84180c75",
2577 => x"ac180c75",
2578 => x"b00c993d",
2579 => x"0d04893d",
2580 => x"70556a54",
2581 => x"558a5299",
2582 => x"3dffbc05",
2583 => x"51ffb7e2",
2584 => x"3fb00877",
2585 => x"53755256",
2586 => x"fecb3fbc",
2587 => x"3f77b008",
2588 => x"0c75b00c",
2589 => x"993d0d04",
2590 => x"fc3d0d81",
2591 => x"5480e3e0",
2592 => x"08883873",
2593 => x"b00c863d",
2594 => x"0d047653",
2595 => x"97b95286",
2596 => x"3dfc0551",
2597 => x"ffb7ab3f",
2598 => x"b008548c",
2599 => x"3f74b008",
2600 => x"0c73b00c",
2601 => x"863d0d04",
2602 => x"80d3f008",
2603 => x"b00c04f7",
2604 => x"3d0d7b80",
2605 => x"d3f00882",
2606 => x"c811085a",
2607 => x"545a7780",
2608 => x"2e80da38",
2609 => x"81881884",
2610 => x"1908ff05",
2611 => x"81712b59",
2612 => x"55598074",
2613 => x"2480ea38",
2614 => x"807424b5",
2615 => x"3873822b",
2616 => x"78118805",
2617 => x"56568180",
2618 => x"19087706",
2619 => x"5372802e",
2620 => x"b6387816",
2621 => x"70085353",
2622 => x"79517408",
2623 => x"53722dff",
2624 => x"14fc17fc",
2625 => x"1779812c",
2626 => x"5a575754",
2627 => x"738025d6",
2628 => x"38770858",
2629 => x"77ffad38",
2630 => x"80d3f008",
2631 => x"53bc1308",
2632 => x"a5387951",
2633 => x"f9dc3f74",
2634 => x"0853722d",
2635 => x"ff14fc17",
2636 => x"fc177981",
2637 => x"2c5a5757",
2638 => x"54738025",
2639 => x"ffa838d1",
2640 => x"398057ff",
2641 => x"93397251",
2642 => x"bc130853",
2643 => x"722d7951",
2644 => x"f9b03fff",
2645 => x"3d0d80e3",
2646 => x"bc0bfc05",
2647 => x"70085252",
2648 => x"70ff2e91",
2649 => x"38702dfc",
2650 => x"12700852",
2651 => x"5270ff2e",
2652 => x"098106f1",
2653 => x"38833d0d",
2654 => x"0404ffb7",
2655 => x"d53f0400",
2656 => x"00ffffff",
2657 => x"ff00ffff",
2658 => x"ffff00ff",
2659 => x"ffffff00",
2660 => x"00000040",
2661 => x"7a707574",
2662 => x"6573740a",
2663 => x"00000000",
2664 => x"48656c6c",
2665 => x"6f20776f",
2666 => x"726c6420",
2667 => x"310a0000",
2668 => x"48656c6c",
2669 => x"6f20776f",
2670 => x"726c6420",
2671 => x"320a0000",
2672 => x"61626f72",
2673 => x"7428290a",
2674 => x"00000000",
2675 => x"0a000000",
2676 => x"43000000",
2677 => x"64756d6d",
2678 => x"792e6578",
2679 => x"65000000",
2680 => x"00000000",
2681 => x"00000000",
2682 => x"00000000",
2683 => x"000031c4",
2684 => x"000029f4",
2685 => x"00000000",
2686 => x"00002c5c",
2687 => x"00002cb8",
2688 => x"00002d14",
2689 => x"00000000",
2690 => x"00000000",
2691 => x"00000000",
2692 => x"00000000",
2693 => x"00000000",
2694 => x"00000000",
2695 => x"00000000",
2696 => x"00000000",
2697 => x"00000000",
2698 => x"000029d0",
2699 => x"00000000",
2700 => x"00000000",
2701 => x"00000000",
2702 => x"00000000",
2703 => x"00000000",
2704 => x"00000000",
2705 => x"00000000",
2706 => x"00000000",
2707 => x"00000000",
2708 => x"00000000",
2709 => x"00000000",
2710 => x"00000000",
2711 => x"00000000",
2712 => x"00000000",
2713 => x"00000000",
2714 => x"00000000",
2715 => x"00000000",
2716 => x"00000000",
2717 => x"00000000",
2718 => x"00000000",
2719 => x"00000000",
2720 => x"00000000",
2721 => x"00000000",
2722 => x"00000000",
2723 => x"00000000",
2724 => x"00000000",
2725 => x"00000000",
2726 => x"00000000",
2727 => x"00000001",
2728 => x"330eabcd",
2729 => x"1234e66d",
2730 => x"deec0005",
2731 => x"000b0000",
2732 => x"00000000",
2733 => x"00000000",
2734 => x"00000000",
2735 => x"00000000",
2736 => x"00000000",
2737 => x"00000000",
2738 => x"00000000",
2739 => x"00000000",
2740 => x"00000000",
2741 => x"00000000",
2742 => x"00000000",
2743 => x"00000000",
2744 => x"00000000",
2745 => x"00000000",
2746 => x"00000000",
2747 => x"00000000",
2748 => x"00000000",
2749 => x"00000000",
2750 => x"00000000",
2751 => x"00000000",
2752 => x"00000000",
2753 => x"00000000",
2754 => x"00000000",
2755 => x"00000000",
2756 => x"00000000",
2757 => x"00000000",
2758 => x"00000000",
2759 => x"00000000",
2760 => x"00000000",
2761 => x"00000000",
2762 => x"00000000",
2763 => x"00000000",
2764 => x"00000000",
2765 => x"00000000",
2766 => x"00000000",
2767 => x"00000000",
2768 => x"00000000",
2769 => x"00000000",
2770 => x"00000000",
2771 => x"00000000",
2772 => x"00000000",
2773 => x"00000000",
2774 => x"00000000",
2775 => x"00000000",
2776 => x"00000000",
2777 => x"00000000",
2778 => x"00000000",
2779 => x"00000000",
2780 => x"00000000",
2781 => x"00000000",
2782 => x"00000000",
2783 => x"00000000",
2784 => x"00000000",
2785 => x"00000000",
2786 => x"00000000",
2787 => x"00000000",
2788 => x"00000000",
2789 => x"00000000",
2790 => x"00000000",
2791 => x"00000000",
2792 => x"00000000",
2793 => x"00000000",
2794 => x"00000000",
2795 => x"00000000",
2796 => x"00000000",
2797 => x"00000000",
2798 => x"00000000",
2799 => x"00000000",
2800 => x"00000000",
2801 => x"00000000",
2802 => x"00000000",
2803 => x"00000000",
2804 => x"00000000",
2805 => x"00000000",
2806 => x"00000000",
2807 => x"00000000",
2808 => x"00000000",
2809 => x"00000000",
2810 => x"00000000",
2811 => x"00000000",
2812 => x"00000000",
2813 => x"00000000",
2814 => x"00000000",
2815 => x"00000000",
2816 => x"00000000",
2817 => x"00000000",
2818 => x"00000000",
2819 => x"00000000",
2820 => x"00000000",
2821 => x"00000000",
2822 => x"00000000",
2823 => x"00000000",
2824 => x"00000000",
2825 => x"00000000",
2826 => x"00000000",
2827 => x"00000000",
2828 => x"00000000",
2829 => x"00000000",
2830 => x"00000000",
2831 => x"00000000",
2832 => x"00000000",
2833 => x"00000000",
2834 => x"00000000",
2835 => x"00000000",
2836 => x"00000000",
2837 => x"00000000",
2838 => x"00000000",
2839 => x"00000000",
2840 => x"00000000",
2841 => x"00000000",
2842 => x"00000000",
2843 => x"00000000",
2844 => x"00000000",
2845 => x"00000000",
2846 => x"00000000",
2847 => x"00000000",
2848 => x"00000000",
2849 => x"00000000",
2850 => x"00000000",
2851 => x"00000000",
2852 => x"00000000",
2853 => x"00000000",
2854 => x"00000000",
2855 => x"00000000",
2856 => x"00000000",
2857 => x"00000000",
2858 => x"00000000",
2859 => x"00000000",
2860 => x"00000000",
2861 => x"00000000",
2862 => x"00000000",
2863 => x"00000000",
2864 => x"00000000",
2865 => x"00000000",
2866 => x"00000000",
2867 => x"00000000",
2868 => x"00000000",
2869 => x"00000000",
2870 => x"00000000",
2871 => x"00000000",
2872 => x"00000000",
2873 => x"00000000",
2874 => x"00000000",
2875 => x"00000000",
2876 => x"00000000",
2877 => x"00000000",
2878 => x"00000000",
2879 => x"00000000",
2880 => x"00000000",
2881 => x"00000000",
2882 => x"00000000",
2883 => x"00000000",
2884 => x"00000000",
2885 => x"00000000",
2886 => x"00000000",
2887 => x"00000000",
2888 => x"00000000",
2889 => x"00000000",
2890 => x"00000000",
2891 => x"00000000",
2892 => x"00000000",
2893 => x"00000000",
2894 => x"00000000",
2895 => x"00000000",
2896 => x"00000000",
2897 => x"00000000",
2898 => x"00000000",
2899 => x"00000000",
2900 => x"00000000",
2901 => x"00000000",
2902 => x"00000000",
2903 => x"00000000",
2904 => x"00000000",
2905 => x"00000000",
2906 => x"00000000",
2907 => x"00000000",
2908 => x"00000000",
2909 => x"00000000",
2910 => x"00000000",
2911 => x"00000000",
2912 => x"00000000",
2913 => x"00000000",
2914 => x"00000000",
2915 => x"00000000",
2916 => x"00000000",
2917 => x"00000000",
2918 => x"00000000",
2919 => x"00000000",
2920 => x"ffffffff",
2921 => x"00000000",
2922 => x"00020000",
2923 => x"00000000",
2924 => x"00000000",
2925 => x"00002dac",
2926 => x"00002dac",
2927 => x"00002db4",
2928 => x"00002db4",
2929 => x"00002dbc",
2930 => x"00002dbc",
2931 => x"00002dc4",
2932 => x"00002dc4",
2933 => x"00002dcc",
2934 => x"00002dcc",
2935 => x"00002dd4",
2936 => x"00002dd4",
2937 => x"00002ddc",
2938 => x"00002ddc",
2939 => x"00002de4",
2940 => x"00002de4",
2941 => x"00002dec",
2942 => x"00002dec",
2943 => x"00002df4",
2944 => x"00002df4",
2945 => x"00002dfc",
2946 => x"00002dfc",
2947 => x"00002e04",
2948 => x"00002e04",
2949 => x"00002e0c",
2950 => x"00002e0c",
2951 => x"00002e14",
2952 => x"00002e14",
2953 => x"00002e1c",
2954 => x"00002e1c",
2955 => x"00002e24",
2956 => x"00002e24",
2957 => x"00002e2c",
2958 => x"00002e2c",
2959 => x"00002e34",
2960 => x"00002e34",
2961 => x"00002e3c",
2962 => x"00002e3c",
2963 => x"00002e44",
2964 => x"00002e44",
2965 => x"00002e4c",
2966 => x"00002e4c",
2967 => x"00002e54",
2968 => x"00002e54",
2969 => x"00002e5c",
2970 => x"00002e5c",
2971 => x"00002e64",
2972 => x"00002e64",
2973 => x"00002e6c",
2974 => x"00002e6c",
2975 => x"00002e74",
2976 => x"00002e74",
2977 => x"00002e7c",
2978 => x"00002e7c",
2979 => x"00002e84",
2980 => x"00002e84",
2981 => x"00002e8c",
2982 => x"00002e8c",
2983 => x"00002e94",
2984 => x"00002e94",
2985 => x"00002e9c",
2986 => x"00002e9c",
2987 => x"00002ea4",
2988 => x"00002ea4",
2989 => x"00002eac",
2990 => x"00002eac",
2991 => x"00002eb4",
2992 => x"00002eb4",
2993 => x"00002ebc",
2994 => x"00002ebc",
2995 => x"00002ec4",
2996 => x"00002ec4",
2997 => x"00002ecc",
2998 => x"00002ecc",
2999 => x"00002ed4",
3000 => x"00002ed4",
3001 => x"00002edc",
3002 => x"00002edc",
3003 => x"00002ee4",
3004 => x"00002ee4",
3005 => x"00002eec",
3006 => x"00002eec",
3007 => x"00002ef4",
3008 => x"00002ef4",
3009 => x"00002efc",
3010 => x"00002efc",
3011 => x"00002f04",
3012 => x"00002f04",
3013 => x"00002f0c",
3014 => x"00002f0c",
3015 => x"00002f14",
3016 => x"00002f14",
3017 => x"00002f1c",
3018 => x"00002f1c",
3019 => x"00002f24",
3020 => x"00002f24",
3021 => x"00002f2c",
3022 => x"00002f2c",
3023 => x"00002f34",
3024 => x"00002f34",
3025 => x"00002f3c",
3026 => x"00002f3c",
3027 => x"00002f44",
3028 => x"00002f44",
3029 => x"00002f4c",
3030 => x"00002f4c",
3031 => x"00002f54",
3032 => x"00002f54",
3033 => x"00002f5c",
3034 => x"00002f5c",
3035 => x"00002f64",
3036 => x"00002f64",
3037 => x"00002f6c",
3038 => x"00002f6c",
3039 => x"00002f74",
3040 => x"00002f74",
3041 => x"00002f7c",
3042 => x"00002f7c",
3043 => x"00002f84",
3044 => x"00002f84",
3045 => x"00002f8c",
3046 => x"00002f8c",
3047 => x"00002f94",
3048 => x"00002f94",
3049 => x"00002f9c",
3050 => x"00002f9c",
3051 => x"00002fa4",
3052 => x"00002fa4",
3053 => x"00002fac",
3054 => x"00002fac",
3055 => x"00002fb4",
3056 => x"00002fb4",
3057 => x"00002fbc",
3058 => x"00002fbc",
3059 => x"00002fc4",
3060 => x"00002fc4",
3061 => x"00002fcc",
3062 => x"00002fcc",
3063 => x"00002fd4",
3064 => x"00002fd4",
3065 => x"00002fdc",
3066 => x"00002fdc",
3067 => x"00002fe4",
3068 => x"00002fe4",
3069 => x"00002fec",
3070 => x"00002fec",
3071 => x"00002ff4",
3072 => x"00002ff4",
3073 => x"00002ffc",
3074 => x"00002ffc",
3075 => x"00003004",
3076 => x"00003004",
3077 => x"0000300c",
3078 => x"0000300c",
3079 => x"00003014",
3080 => x"00003014",
3081 => x"0000301c",
3082 => x"0000301c",
3083 => x"00003024",
3084 => x"00003024",
3085 => x"0000302c",
3086 => x"0000302c",
3087 => x"00003034",
3088 => x"00003034",
3089 => x"0000303c",
3090 => x"0000303c",
3091 => x"00003044",
3092 => x"00003044",
3093 => x"0000304c",
3094 => x"0000304c",
3095 => x"00003054",
3096 => x"00003054",
3097 => x"0000305c",
3098 => x"0000305c",
3099 => x"00003064",
3100 => x"00003064",
3101 => x"0000306c",
3102 => x"0000306c",
3103 => x"00003074",
3104 => x"00003074",
3105 => x"0000307c",
3106 => x"0000307c",
3107 => x"00003084",
3108 => x"00003084",
3109 => x"0000308c",
3110 => x"0000308c",
3111 => x"00003094",
3112 => x"00003094",
3113 => x"0000309c",
3114 => x"0000309c",
3115 => x"000030a4",
3116 => x"000030a4",
3117 => x"000030ac",
3118 => x"000030ac",
3119 => x"000030b4",
3120 => x"000030b4",
3121 => x"000030bc",
3122 => x"000030bc",
3123 => x"000030c4",
3124 => x"000030c4",
3125 => x"000030cc",
3126 => x"000030cc",
3127 => x"000030d4",
3128 => x"000030d4",
3129 => x"000030dc",
3130 => x"000030dc",
3131 => x"000030e4",
3132 => x"000030e4",
3133 => x"000030ec",
3134 => x"000030ec",
3135 => x"000030f4",
3136 => x"000030f4",
3137 => x"000030fc",
3138 => x"000030fc",
3139 => x"00003104",
3140 => x"00003104",
3141 => x"0000310c",
3142 => x"0000310c",
3143 => x"00003114",
3144 => x"00003114",
3145 => x"0000311c",
3146 => x"0000311c",
3147 => x"00003124",
3148 => x"00003124",
3149 => x"0000312c",
3150 => x"0000312c",
3151 => x"00003134",
3152 => x"00003134",
3153 => x"0000313c",
3154 => x"0000313c",
3155 => x"00003144",
3156 => x"00003144",
3157 => x"0000314c",
3158 => x"0000314c",
3159 => x"00003154",
3160 => x"00003154",
3161 => x"0000315c",
3162 => x"0000315c",
3163 => x"00003164",
3164 => x"00003164",
3165 => x"0000316c",
3166 => x"0000316c",
3167 => x"00003174",
3168 => x"00003174",
3169 => x"0000317c",
3170 => x"0000317c",
3171 => x"00003184",
3172 => x"00003184",
3173 => x"0000318c",
3174 => x"0000318c",
3175 => x"00003194",
3176 => x"00003194",
3177 => x"0000319c",
3178 => x"0000319c",
3179 => x"000031a4",
3180 => x"000031a4",
3181 => x"000029d4",
3182 => x"ffffffff",
3183 => x"00000000",
3184 => x"ffffffff",
3185 => x"00000000",


others => x"00000000"
);
begin
   do_port_a:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         if (a_we_i='1') and (b_we_i='1') and (a_addr_i=b_addr_i) and (a_write_i/=b_write_i) then
            report "DualPortRAM write collision" severity failure;
         end if;
         iaddr:=to_integer(a_addr_i);
         if a_we_i='1' then
            ram(iaddr):=a_write_i;
            -- Write First mode
            a_read_o <= a_write_i;
         else
            a_read_o <= ram(iaddr);
         end if;
      end if;
   end process do_port_a;

   do_port_b:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         iaddr:=to_integer(b_addr_i);
         if b_we_i='1' then
            ram(iaddr):=b_write_i;
            b_read_o <= b_write_i;
         else
            b_read_o <= ram(iaddr);
         end if;
      end if;
   end process do_port_b;
end architecture Xilinx; -- Entity: DualPortRAM
